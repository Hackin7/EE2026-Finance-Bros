module video(
    // Control
    input reset, input clk,
    // LEDs, Switches, Buttons
    input btnU, btnL, btnR, btnD, input [15:0] sw, output [15:0] led,
    // 7 Segment Display
    output [6:0] seg, output dp, output [3:0] an,
    // OLED
    inout [7:0] JB,
    output hsync,
    output vsync,
    output [11:0] rgb
);
    //// OLED Setup ////////////////////////////////////////////////////////
    wire [7:0] Jb;
    assign JB[7:0] = Jb;
    wire clk_6_25mhz;
    clk_counter #(16, 5) clk6p25m (clk, clk_6_25mhz);
    reg [15:0] frame_memory [0:7679]; // Adjust size based on image dimensions (96x64 for example)
    
    reg [6:0] frame_counter = 0;
    reg [31:0] frame_timer = 0;
    
    always @(posedge clk) begin
        if (reset) begin
            frame_counter <= 0;
            frame_timer <= 0;
        end else begin
            if (btnU) begin
                if (frame_timer >= 20_000_000) begin // 5 FPS (100 MHz / 5 = 20,000,000)
                    frame_timer <= 0;
                    if (frame_counter < 74) begin
                        frame_counter <= frame_counter + 1;
                    end else begin
                        frame_counter <= 0;
                    end
                end else begin
                    frame_timer <= frame_timer + 1;
                end
            end
        end
    end
    
    // Load frame data based on frame counter
    always @(posedge clk) begin
        case (frame_counter)
            // Frame loading statements will be generated by the Python script
            0: $readmemh("frame_0000.mem", frame_memory);
1: $readmemh("frame_0001.mem", frame_memory);
2: $readmemh("frame_0002.mem", frame_memory);
3: $readmemh("frame_0003.mem", frame_memory);
4: $readmemh("frame_0004.mem", frame_memory);
5: $readmemh("frame_0005.mem", frame_memory);
6: $readmemh("frame_0006.mem", frame_memory);
7: $readmemh("frame_0007.mem", frame_memory);
8: $readmemh("frame_0008.mem", frame_memory);
9: $readmemh("frame_0009.mem", frame_memory);
10: $readmemh("frame_0010.mem", frame_memory);
11: $readmemh("frame_0011.mem", frame_memory);
12: $readmemh("frame_0012.mem", frame_memory);
13: $readmemh("frame_0013.mem", frame_memory);
14: $readmemh("frame_0014.mem", frame_memory);
15: $readmemh("frame_0015.mem", frame_memory);
16: $readmemh("frame_0016.mem", frame_memory);
17: $readmemh("frame_0017.mem", frame_memory);
18: $readmemh("frame_0018.mem", frame_memory);
19: $readmemh("frame_0019.mem", frame_memory);
20: $readmemh("frame_0020.mem", frame_memory);
21: $readmemh("frame_0021.mem", frame_memory);
22: $readmemh("frame_0022.mem", frame_memory);
23: $readmemh("frame_0023.mem", frame_memory);
24: $readmemh("frame_0024.mem", frame_memory);
25: $readmemh("frame_0025.mem", frame_memory);
26: $readmemh("frame_0026.mem", frame_memory);
27: $readmemh("frame_0027.mem", frame_memory);
28: $readmemh("frame_0028.mem", frame_memory);
29: $readmemh("frame_0029.mem", frame_memory);
30: $readmemh("frame_0030.mem", frame_memory);
31: $readmemh("frame_0031.mem", frame_memory);
32: $readmemh("frame_0032.mem", frame_memory);
33: $readmemh("frame_0033.mem", frame_memory);
34: $readmemh("frame_0034.mem", frame_memory);
35: $readmemh("frame_0035.mem", frame_memory);
36: $readmemh("frame_0036.mem", frame_memory);
37: $readmemh("frame_0037.mem", frame_memory);
38: $readmemh("frame_0038.mem", frame_memory);
39: $readmemh("frame_0039.mem", frame_memory);
40: $readmemh("frame_0040.mem", frame_memory);
41: $readmemh("frame_0041.mem", frame_memory);
42: $readmemh("frame_0042.mem", frame_memory);
43: $readmemh("frame_0043.mem", frame_memory);
44: $readmemh("frame_0044.mem", frame_memory);
45: $readmemh("frame_0045.mem", frame_memory);
46: $readmemh("frame_0046.mem", frame_memory);
47: $readmemh("frame_0047.mem", frame_memory);
48: $readmemh("frame_0048.mem", frame_memory);
49: $readmemh("frame_0049.mem", frame_memory);
50: $readmemh("frame_0050.mem", frame_memory);
51: $readmemh("frame_0051.mem", frame_memory);
52: $readmemh("frame_0052.mem", frame_memory);
53: $readmemh("frame_0053.mem", frame_memory);
54: $readmemh("frame_0054.mem", frame_memory);
55: $readmemh("frame_0055.mem", frame_memory);
56: $readmemh("frame_0056.mem", frame_memory);
57: $readmemh("frame_0057.mem", frame_memory);
58: $readmemh("frame_0058.mem", frame_memory);
59: $readmemh("frame_0059.mem", frame_memory);
60: $readmemh("frame_0060.mem", frame_memory);
61: $readmemh("frame_0061.mem", frame_memory);
62: $readmemh("frame_0062.mem", frame_memory);
63: $readmemh("frame_0063.mem", frame_memory);
64: $readmemh("frame_0064.mem", frame_memory);
65: $readmemh("frame_0065.mem", frame_memory);
66: $readmemh("frame_0066.mem", frame_memory);
67: $readmemh("frame_0067.mem", frame_memory);
68: $readmemh("frame_0068.mem", frame_memory);
69: $readmemh("frame_0069.mem", frame_memory);
70: $readmemh("frame_0070.mem", frame_memory);
71: $readmemh("frame_0071.mem", frame_memory);
72: $readmemh("frame_0072.mem", frame_memory);
73: $readmemh("frame_0073.mem", frame_memory);
74: $readmemh("frame_0074.mem", frame_memory);

        endcase
    end
    
    wire [12:0] oled_pixel_index;
    wire [15:0] pixel_data;
    
    assign pixel_data = frame_memory[oled_pixel_index];
    
    vga_oled_adaptor adaptor(
        .clk(clk),
        .reset(reset),
        .JB(JB),
        .pixel_index(oled_pixel_index),
        .pixel_data(pixel_data),
        .hsync(hsync),
        .vsync(vsync),
        .rgb(rgb)
    );
endmodule