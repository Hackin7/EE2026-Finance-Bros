module video(
    // Control
    input reset, input clk,
    // LEDs, Switches, Buttons
    input btnU, btnL, btnR, btnD, input [15:0] sw, output [15:0] led,
    // 7 Segment Display
    output [6:0] seg, output dp, output [3:0] an,
    // OLED
    inout [7:0] JB,
    output hsync,
    output vsync,
    output [11:0] rgb
);
    //// OLED Setup ////////////////////////////////////////////////////////
    wire [7:0] Jb;
    assign JB[7:0] = Jb;
    wire clk_6_25mhz;
    clk_counter #(16, 5) clk6p25m (clk, clk_6_25mhz);
    reg [15:0] frame_memory [0:7679]; // Adjust size based on image dimensions (96x64 for example)
    
    reg [6:0] frame_counter = 0;
    reg [31:0] frame_timer = 0;
    
    always @(posedge clk) begin
        if (reset) begin
            frame_counter <= 0;
            frame_timer <= 0;
        end else begin
            if (btnU) begin
                if (frame_timer >= 20_000_000) begin // 5 FPS (100 MHz / 5 = 20,000,000)
                    frame_timer <= 0;
                    if (frame_counter < 74) begin
                        frame_counter <= frame_counter + 1;
                    end else begin
                        frame_counter <= 0;
                    end
                end else begin
                    frame_timer <= frame_timer + 1;
                end
            end
        end
    end
    
    // Load frame data based on frame counter
    always @(posedge clk) begin
        case (frame_counter)
            // Frame loading statements will be generated by the Python script
            {{FRAME_LOADING_STATEMENTS}}
        endcase
    end
    
    wire [12:0] oled_pixel_index;
    wire [15:0] pixel_data;
    
    assign pixel_data = frame_memory[oled_pixel_index];
    
    vga_oled_adaptor adaptor(
        .clk(clk),
        .reset(reset),
        .JB(JB),
        .pixel_index(oled_pixel_index),
        .pixel_data(pixel_data),
        .hsync(hsync),
        .vsync(vsync),
        .rgb(rgb)
    );
endmodule